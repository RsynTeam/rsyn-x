VERSION 5.7 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS	2000 ;
END UNITS

MANUFACTURINGGRID	0.0025 ;

SITE core
  SIZE 0.19 BY 1.71 ;
  CLASS CORE ;
END core

LAYER metal1
  TYPE			ROUTING ;
  DIRECTION		HORIZONTAL ;
  PITCH			0.200 ;
  OFFSET		0.000 ;
  WIDTH			0.100 ;
END metal1

LAYER metal2
  TYPE			ROUTING ;
  DIRECTION		VERTICAL ;
  PITCH			0.200 ;
  OFFSET		0.100 ;
  WIDTH			0.1 ;
END metal2

LAYER metal3
  TYPE			ROUTING ;
  DIRECTION		HORIZONTAL ;
  PITCH			0.200 ;
  OFFSET		0.000 ;
  WIDTH			0.1 ;
END metal3

MACRO INV_X1
    CLASS CORE ;
    FOREIGN INV_X1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.760 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.150 0.53 1.255 ;
        RECT 0.415 0.150 0.61 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.340 0.34 0.405 ;
        END
    END a
END INV_X1

MACRO INV_X2
    CLASS CORE ;
    FOREIGN INV_X2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.150 1.12 1.255 ;
        RECT 0.835 0.150 1.225 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.340 0.68 0.405 ;
        END
    END a
END INV_X2

MACRO INV_X3
    CLASS CORE ;
    FOREIGN INV_X3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.900 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.150 1.355 1.255 ;
        RECT 1.040 0.150 1.495 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.340 0.85 0.405 ;
        END
    END a
END INV_X3

MACRO INV_X4
    CLASS CORE ;
    FOREIGN INV_X4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.900 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.150 1.355 1.255 ;
        RECT 1.040 0.150 1.495 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.340 0.85 0.405 ;
        END
    END a
END INV_X4

MACRO INV_X6
    CLASS CORE ;
    FOREIGN INV_X6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.280 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.150 1.65 1.255 ;
        RECT 1.250 0.150 1.77 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.340 1.02 0.405 ;
        END
    END a
END INV_X6

MACRO INV_X8
    CLASS CORE ;
    FOREIGN INV_X8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.150 1.945 1.255 ;
        RECT 1.460 0.150 2.11 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.340 1.19 0.405 ;
        END
    END a
END INV_X8

MACRO INV_X10
    CLASS CORE ;
    FOREIGN INV_X10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.150 1.945 1.255 ;
        RECT 1.460 0.150 2.11 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.340 1.19 0.405 ;
        END
    END a
END INV_X10

MACRO INV_X20
    CLASS CORE ;
    FOREIGN INV_X20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.315 0.150 2.77 1.255 ;
        RECT 2.085 0.150 2.995 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.050 0.340 1.7 0.405 ;
        END
    END a
END INV_X20

MACRO INV_X40
    CLASS CORE ;
    FOREIGN INV_X40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.010 0.150 3.595 1.255 ;
        RECT 2.710 0.150 3.88 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.365 0.340 2.21 0.405 ;
        END
    END a
END INV_X40

MACRO INV_X80
    CLASS CORE ;
    FOREIGN INV_X80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.840 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.170 0.150 4.95 1.255 ;
        RECT 3.750 0.150 5.375 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.890 0.340 3.06 0.405 ;
        END
    END a
END INV_X80

MACRO INV_Y1
    CLASS CORE ;
    FOREIGN INV_Y1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.760 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.150 0.53 1.255 ;
        RECT 0.415 0.150 0.61 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.340 0.34 0.405 ;
        END
    END a
END INV_Y1

MACRO INV_Y2
    CLASS CORE ;
    FOREIGN INV_Y2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.150 1.12 1.255 ;
        RECT 0.835 0.150 1.225 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.340 0.68 0.405 ;
        END
    END a
END INV_Y2

MACRO INV_Y3
    CLASS CORE ;
    FOREIGN INV_Y3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.900 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.150 1.355 1.255 ;
        RECT 1.040 0.150 1.495 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.340 0.85 0.405 ;
        END
    END a
END INV_Y3

MACRO INV_Y4
    CLASS CORE ;
    FOREIGN INV_Y4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.900 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.150 1.355 1.255 ;
        RECT 1.040 0.150 1.495 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.340 0.85 0.405 ;
        END
    END a
END INV_Y4

MACRO INV_Y6
    CLASS CORE ;
    FOREIGN INV_Y6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.280 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.150 1.65 1.255 ;
        RECT 1.250 0.150 1.77 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.340 1.02 0.405 ;
        END
    END a
END INV_Y6

MACRO INV_Y8
    CLASS CORE ;
    FOREIGN INV_Y8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.150 1.945 1.255 ;
        RECT 1.460 0.150 2.11 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.340 1.19 0.405 ;
        END
    END a
END INV_Y8

MACRO INV_Y10
    CLASS CORE ;
    FOREIGN INV_Y10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.150 1.945 1.255 ;
        RECT 1.460 0.150 2.11 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.340 1.19 0.405 ;
        END
    END a
END INV_Y10

MACRO INV_Y20
    CLASS CORE ;
    FOREIGN INV_Y20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.315 0.150 2.77 1.255 ;
        RECT 2.085 0.150 2.995 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.050 0.340 1.7 0.405 ;
        END
    END a
END INV_Y20

MACRO INV_Y40
    CLASS CORE ;
    FOREIGN INV_Y40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.010 0.150 3.595 1.255 ;
        RECT 2.710 0.150 3.88 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.365 0.340 2.21 0.405 ;
        END
    END a
END INV_Y40

MACRO INV_Y80
    CLASS CORE ;
    FOREIGN INV_Y80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.840 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.170 0.150 4.95 1.255 ;
        RECT 3.750 0.150 5.375 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.890 0.340 3.06 0.405 ;
        END
    END a
END INV_Y80

MACRO INV_Z1
    CLASS CORE ;
    FOREIGN INV_Z1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 0.760 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.150 0.53 1.255 ;
        RECT 0.415 0.150 0.61 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.340 0.34 0.405 ;
        END
    END a
END INV_Z1

MACRO INV_Z2
    CLASS CORE ;
    FOREIGN INV_Z2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.150 1.12 1.255 ;
        RECT 0.835 0.150 1.225 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.340 0.68 0.405 ;
        END
    END a
END INV_Z2

MACRO INV_Z3
    CLASS CORE ;
    FOREIGN INV_Z3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.900 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.150 1.355 1.255 ;
        RECT 1.040 0.150 1.495 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.340 0.85 0.405 ;
        END
    END a
END INV_Z3

MACRO INV_Z4
    CLASS CORE ;
    FOREIGN INV_Z4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.900 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.150 1.355 1.255 ;
        RECT 1.040 0.150 1.495 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.340 0.85 0.405 ;
        END
    END a
END INV_Z4

MACRO INV_Z6
    CLASS CORE ;
    FOREIGN INV_Z6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.280 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.150 1.65 1.255 ;
        RECT 1.250 0.150 1.77 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.340 1.02 0.405 ;
        END
    END a
END INV_Z6

MACRO INV_Z8
    CLASS CORE ;
    FOREIGN INV_Z8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.150 1.945 1.255 ;
        RECT 1.460 0.150 2.11 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.340 1.19 0.405 ;
        END
    END a
END INV_Z8

MACRO INV_Z10
    CLASS CORE ;
    FOREIGN INV_Z10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.150 1.945 1.255 ;
        RECT 1.460 0.150 2.11 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.340 1.19 0.405 ;
        END
    END a
END INV_Z10

MACRO INV_Z20
    CLASS CORE ;
    FOREIGN INV_Z20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.315 0.150 2.77 1.255 ;
        RECT 2.085 0.150 2.995 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.050 0.340 1.7 0.405 ;
        END
    END a
END INV_Z20

MACRO INV_Z40
    CLASS CORE ;
    FOREIGN INV_Z40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.010 0.150 3.595 1.255 ;
        RECT 2.710 0.150 3.88 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.365 0.340 2.21 0.405 ;
        END
    END a
END INV_Z40

MACRO INV_Z80
    CLASS CORE ;
    FOREIGN INV_Z80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.840 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.170 0.150 4.95 1.255 ;
        RECT 3.750 0.150 5.375 0.28 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.890 0.340 3.06 0.405 ;
        END
    END a
END INV_Z80

MACRO NAND2_X1
    CLASS CORE ;
    FOREIGN NAND2_X1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.450 0.110 0.58 1.215 ;
        RECT 0.430 0.725 0.625 1.245 ;
        RECT 0.450 0.110 0.905 0.175 ;
        RECT 0.805 0.110 0.935 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.070 0.535 0.33 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.645 0.540 0.905 0.67 ;
        END
    END b
END NAND2_X1

MACRO NAND2_X2
    CLASS CORE ;
    FOREIGN NAND2_X2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.050 0.110 1.31 1.215 ;
        RECT 1.000 0.725 1.455 1.245 ;
        RECT 1.050 0.110 2.09 0.175 ;
        RECT 1.875 0.110 2.135 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.160 0.535 0.81 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.505 0.540 2.09 0.67 ;
        END
    END b
END NAND2_X2

MACRO NAND2_X3
    CLASS CORE ;
    FOREIGN NAND2_X3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.350 0.110 1.675 1.215 ;
        RECT 1.285 0.725 1.87 1.245 ;
        RECT 1.350 0.110 2.715 0.175 ;
        RECT 2.410 0.110 2.735 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.205 0.535 1.05 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.935 0.540 2.715 0.67 ;
        END
    END b
END NAND2_X3

MACRO NAND2_X4
    CLASS CORE ;
    FOREIGN NAND2_X4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.500 0.110 1.825 1.215 ;
        RECT 1.425 0.725 2.075 1.245 ;
        RECT 1.500 0.110 2.995 0.175 ;
        RECT 2.675 0.110 3.0 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.225 0.535 1.2 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.540 2.995 0.67 ;
        END
    END b
END NAND2_X4

MACRO NAND2_X6
    CLASS CORE ;
    FOREIGN NAND2_X6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.800 0.110 2.19 1.215 ;
        RECT 1.710 0.725 2.49 1.245 ;
        RECT 1.800 0.110 3.62 0.175 ;
        RECT 3.210 0.110 3.6 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.270 0.535 1.44 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.540 3.62 0.67 ;
        END
    END b
END NAND2_X6

MACRO NAND2_X8
    CLASS CORE ;
    FOREIGN NAND2_X8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.950 0.110 2.405 1.215 ;
        RECT 1.855 0.725 2.7 1.245 ;
        RECT 1.950 0.110 3.9 0.175 ;
        RECT 3.480 0.110 3.935 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.290 0.535 1.525 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.795 0.540 3.9 0.67 ;
        END
    END b
END NAND2_X8

MACRO NAND2_X10
    CLASS CORE ;
    FOREIGN NAND2_X10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.250 0.110 2.77 1.215 ;
        RECT 2.140 0.725 3.18 1.245 ;
        RECT 2.250 0.110 4.525 0.175 ;
        RECT 4.015 0.110 4.535 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.340 0.535 1.77 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.225 0.540 4.525 0.67 ;
        END
    END b
END NAND2_X10

MACRO NAND2_X20
    CLASS CORE ;
    FOREIGN NAND2_X20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.000 0.110 3.65 1.215 ;
        RECT 2.850 0.725 4.215 1.245 ;
        RECT 3.000 0.110 5.99 0.175 ;
        RECT 5.350 0.110 6.0 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.450 0.535 2.335 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.540 6.055 0.67 ;
        END
    END b
END NAND2_X20

MACRO NAND2_X40
    CLASS CORE ;
    FOREIGN NAND2_X40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.200 0.110 5.11 1.215 ;
        RECT 3.990 0.725 5.875 1.245 ;
        RECT 4.200 0.110 8.425 0.175 ;
        RECT 7.490 0.110 8.4 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.535 3.295 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.020 0.540 8.425 0.67 ;
        END
    END b
END NAND2_X40

MACRO NAND2_X80
    CLASS CORE ;
    FOREIGN NAND2_X80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.700 0.110 6.935 1.215 ;
        RECT 5.415 0.725 7.95 1.245 ;
        RECT 5.700 0.110 11.42 0.175 ;
        RECT 10.165 0.110 11.4 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.855 0.535 4.495 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.170 0.540 11.42 0.67 ;
        END
    END b
END NAND2_X80

MACRO NAND2_Y01
    CLASS CORE ;
    FOREIGN NAND2_Y01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.450 0.110 0.58 1.215 ;
        RECT 0.430 0.725 0.625 1.245 ;
        RECT 0.450 0.110 0.905 0.175 ;
        RECT 0.805 0.110 0.935 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.070 0.535 0.33 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.645 0.540 0.905 0.67 ;
        END
    END b
END NAND2_Y01

MACRO NAND2_Y02
    CLASS CORE ;
    FOREIGN NAND2_Y02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.050 0.110 1.31 1.215 ;
        RECT 1.000 0.725 1.455 1.245 ;
        RECT 1.050 0.110 2.09 0.175 ;
        RECT 1.875 0.110 2.135 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.160 0.535 0.81 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.505 0.540 2.09 0.67 ;
        END
    END b
END NAND2_Y02

MACRO NAND2_Y03
    CLASS CORE ;
    FOREIGN NAND2_Y03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.350 0.110 1.675 1.215 ;
        RECT 1.285 0.725 1.87 1.245 ;
        RECT 1.350 0.110 2.715 0.175 ;
        RECT 2.410 0.110 2.735 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.205 0.535 1.05 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.935 0.540 2.715 0.67 ;
        END
    END b
END NAND2_Y03

MACRO NAND2_Y04
    CLASS CORE ;
    FOREIGN NAND2_Y04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.500 0.110 1.825 1.215 ;
        RECT 1.425 0.725 2.075 1.245 ;
        RECT 1.500 0.110 2.995 0.175 ;
        RECT 2.675 0.110 3.0 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.225 0.535 1.2 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.540 2.995 0.67 ;
        END
    END b
END NAND2_Y04

MACRO NAND2_Y06
    CLASS CORE ;
    FOREIGN NAND2_Y06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.800 0.110 2.19 1.215 ;
        RECT 1.710 0.725 2.49 1.245 ;
        RECT 1.800 0.110 3.62 0.175 ;
        RECT 3.210 0.110 3.6 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.270 0.535 1.44 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.540 3.62 0.67 ;
        END
    END b
END NAND2_Y06

MACRO NAND2_Y08
    CLASS CORE ;
    FOREIGN NAND2_Y08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.950 0.110 2.405 1.215 ;
        RECT 1.855 0.725 2.7 1.245 ;
        RECT 1.950 0.110 3.9 0.175 ;
        RECT 3.480 0.110 3.935 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.290 0.535 1.525 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.795 0.540 3.9 0.67 ;
        END
    END b
END NAND2_Y08

MACRO NAND2_Y10
    CLASS CORE ;
    FOREIGN NAND2_Y10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.250 0.110 2.77 1.215 ;
        RECT 2.140 0.725 3.18 1.245 ;
        RECT 2.250 0.110 4.525 0.175 ;
        RECT 4.015 0.110 4.535 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.340 0.535 1.77 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.225 0.540 4.525 0.67 ;
        END
    END b
END NAND2_Y10

MACRO NAND2_Y20
    CLASS CORE ;
    FOREIGN NAND2_Y20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.000 0.110 3.65 1.215 ;
        RECT 2.850 0.725 4.215 1.245 ;
        RECT 3.000 0.110 5.99 0.175 ;
        RECT 5.350 0.110 6.0 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.450 0.535 2.335 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.540 6.055 0.67 ;
        END
    END b
END NAND2_Y20

MACRO NAND2_Y40
    CLASS CORE ;
    FOREIGN NAND2_Y40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.200 0.110 5.11 1.215 ;
        RECT 3.990 0.725 5.875 1.245 ;
        RECT 4.200 0.110 8.425 0.175 ;
        RECT 7.490 0.110 8.4 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.535 3.295 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.020 0.540 8.425 0.67 ;
        END
    END b
END NAND2_Y40

MACRO NAND2_Y80
    CLASS CORE ;
    FOREIGN NAND2_Y80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.700 0.110 6.935 1.215 ;
        RECT 5.415 0.725 7.95 1.245 ;
        RECT 5.700 0.110 11.42 0.175 ;
        RECT 10.165 0.110 11.4 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.855 0.535 4.495 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.170 0.540 11.42 0.67 ;
        END
    END b
END NAND2_Y80

MACRO NAND2_Z01
    CLASS CORE ;
    FOREIGN NAND2_Z01 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.450 0.110 0.58 1.215 ;
        RECT 0.430 0.725 0.625 1.245 ;
        RECT 0.450 0.110 0.905 0.175 ;
        RECT 0.805 0.110 0.935 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.070 0.535 0.33 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.645 0.540 0.905 0.67 ;
        END
    END b
END NAND2_Z01

MACRO NAND2_Z02
    CLASS CORE ;
    FOREIGN NAND2_Z02 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.050 0.110 1.31 1.215 ;
        RECT 1.000 0.725 1.455 1.245 ;
        RECT 1.050 0.110 2.09 0.175 ;
        RECT 1.875 0.110 2.135 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.160 0.535 0.81 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.505 0.540 2.09 0.67 ;
        END
    END b
END NAND2_Z02

MACRO NAND2_Z03
    CLASS CORE ;
    FOREIGN NAND2_Z03 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.350 0.110 1.675 1.215 ;
        RECT 1.285 0.725 1.87 1.245 ;
        RECT 1.350 0.110 2.715 0.175 ;
        RECT 2.410 0.110 2.735 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.205 0.535 1.05 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.935 0.540 2.715 0.67 ;
        END
    END b
END NAND2_Z03

MACRO NAND2_Z04
    CLASS CORE ;
    FOREIGN NAND2_Z04 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.500 0.110 1.825 1.215 ;
        RECT 1.425 0.725 2.075 1.245 ;
        RECT 1.500 0.110 2.995 0.175 ;
        RECT 2.675 0.110 3.0 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.225 0.535 1.2 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.540 2.995 0.67 ;
        END
    END b
END NAND2_Z04

MACRO NAND2_Z06
    CLASS CORE ;
    FOREIGN NAND2_Z06 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.800 0.110 2.19 1.215 ;
        RECT 1.710 0.725 2.49 1.245 ;
        RECT 1.800 0.110 3.62 0.175 ;
        RECT 3.210 0.110 3.6 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.270 0.535 1.44 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.540 3.62 0.67 ;
        END
    END b
END NAND2_Z06

MACRO NAND2_Z08
    CLASS CORE ;
    FOREIGN NAND2_Z08 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.950 0.110 2.405 1.215 ;
        RECT 1.855 0.725 2.7 1.245 ;
        RECT 1.950 0.110 3.9 0.175 ;
        RECT 3.480 0.110 3.935 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.290 0.535 1.525 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.795 0.540 3.9 0.67 ;
        END
    END b
END NAND2_Z08

MACRO NAND2_Z10
    CLASS CORE ;
    FOREIGN NAND2_Z10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.250 0.110 2.77 1.215 ;
        RECT 2.140 0.725 3.18 1.245 ;
        RECT 2.250 0.110 4.525 0.175 ;
        RECT 4.015 0.110 4.535 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.340 0.535 1.77 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.225 0.540 4.525 0.67 ;
        END
    END b
END NAND2_Z10

MACRO NAND2_Z20
    CLASS CORE ;
    FOREIGN NAND2_Z20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.000 0.110 3.65 1.215 ;
        RECT 2.850 0.725 4.215 1.245 ;
        RECT 3.000 0.110 5.99 0.175 ;
        RECT 5.350 0.110 6.0 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.450 0.535 2.335 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.540 6.055 0.67 ;
        END
    END b
END NAND2_Z20

MACRO NAND2_Z40
    CLASS CORE ;
    FOREIGN NAND2_Z40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.200 0.110 5.11 1.215 ;
        RECT 3.990 0.725 5.875 1.245 ;
        RECT 4.200 0.110 8.425 0.175 ;
        RECT 7.490 0.110 8.4 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.535 3.295 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.020 0.540 8.425 0.67 ;
        END
    END b
END NAND2_Z40

MACRO NAND2_Z80
    CLASS CORE ;
    FOREIGN NAND2_Z80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.700 0.110 6.935 1.215 ;
        RECT 5.415 0.725 7.95 1.245 ;
        RECT 5.700 0.110 11.42 0.175 ;
        RECT 10.165 0.110 11.4 0.5 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.855 0.535 4.495 0.665 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.170 0.540 11.42 0.67 ;
        END
    END b
END NAND2_Z80

MACRO NAND3_X1
    CLASS CORE ;
    FOREIGN NAND3_X1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.415 0.805 0.48 1.26 ;
        RECT 0.415 0.805 0.935 0.87 ;
        RECT 0.875 0.090 0.94 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.040 0.630 0.3 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.350 0.090 0.545 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.640 0.090 0.77 0.74 ;
        END
    END c
END NAND3_X1

MACRO NAND3_X2
    CLASS CORE ;
    FOREIGN NAND3_X2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.975 0.805 1.17 1.26 ;
        RECT 0.975 0.805 2.21 0.87 ;
        RECT 2.035 0.090 2.23 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.090 0.630 0.61 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.820 0.090 1.34 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.490 0.090 1.815 0.74 ;
        END
    END c
END NAND3_X2

MACRO NAND3_X3
    CLASS CORE ;
    FOREIGN NAND3_X3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.250 0.805 1.51 1.26 ;
        RECT 1.250 0.805 2.875 0.87 ;
        RECT 2.620 0.090 2.88 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.115 0.630 0.83 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.055 0.090 1.705 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.915 0.090 2.37 0.74 ;
        END
    END c
END NAND3_X3

MACRO NAND3_X4
    CLASS CORE ;
    FOREIGN NAND3_X4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.805 1.65 1.26 ;
        RECT 1.390 0.805 3.145 0.87 ;
        RECT 2.910 0.090 3.17 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.130 0.630 0.91 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.170 0.090 1.885 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.130 0.090 2.65 0.74 ;
        END
    END c
END NAND3_X4

MACRO NAND3_X6
    CLASS CORE ;
    FOREIGN NAND3_X6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.805 1.995 1.26 ;
        RECT 1.670 0.805 3.815 0.87 ;
        RECT 3.490 0.090 3.815 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.155 0.630 1.065 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.405 0.090 2.25 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.555 0.090 3.14 0.74 ;
        END
    END c
END NAND3_X6

MACRO NAND3_X8
    CLASS CORE ;
    FOREIGN NAND3_X8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.805 0.805 2.13 1.26 ;
        RECT 1.805 0.805 4.145 0.87 ;
        RECT 3.785 0.090 4.11 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.170 0.630 1.145 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.520 0.090 2.43 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.770 0.090 3.42 0.74 ;
        END
    END c
END NAND3_X8

MACRO NAND3_X10
    CLASS CORE ;
    FOREIGN NAND3_X10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.805 2.475 1.26 ;
        RECT 2.085 0.805 4.75 0.87 ;
        RECT 4.365 0.090 4.755 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.195 0.630 1.365 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.755 0.090 2.795 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.195 0.090 3.975 0.74 ;
        END
    END c
END NAND3_X10

MACRO NAND3_X20
    CLASS CORE ;
    FOREIGN NAND3_X20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.805 3.3 1.26 ;
        RECT 2.780 0.805 6.355 0.87 ;
        RECT 5.820 0.090 6.34 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.260 0.630 1.755 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.340 0.090 3.77 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.260 0.090 5.235 0.74 ;
        END
    END c
END NAND3_X20

MACRO NAND3_X40
    CLASS CORE ;
    FOREIGN NAND3_X40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.890 0.805 4.605 1.26 ;
        RECT 3.890 0.805 8.895 0.87 ;
        RECT 8.150 0.090 8.865 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.365 0.630 2.51 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.275 0.090 5.225 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.965 0.090 7.395 0.74 ;
        END
    END c
END NAND3_X40

MACRO NAND3_X80
    CLASS CORE ;
    FOREIGN NAND3_X80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.280 0.805 6.255 1.26 ;
        RECT 5.280 0.805 12.04 0.87 ;
        RECT 11.060 0.090 12.035 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.495 0.630 3.355 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.445 0.090 7.11 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.095 0.090 9.98 0.74 ;
        END
    END c
END NAND3_X80

MACRO NAND3_Y1
    CLASS CORE ;
    FOREIGN NAND3_Y1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.415 0.805 0.48 1.26 ;
        RECT 0.415 0.805 0.935 0.87 ;
        RECT 0.875 0.090 0.94 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.040 0.630 0.3 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.350 0.090 0.545 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.640 0.090 0.77 0.74 ;
        END
    END c
END NAND3_Y1

MACRO NAND3_Y2
    CLASS CORE ;
    FOREIGN NAND3_Y2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.975 0.805 1.17 1.26 ;
        RECT 0.975 0.805 2.21 0.87 ;
        RECT 2.035 0.090 2.23 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.090 0.630 0.61 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.820 0.090 1.34 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.490 0.090 1.815 0.74 ;
        END
    END c
END NAND3_Y2

MACRO NAND3_Y3
    CLASS CORE ;
    FOREIGN NAND3_Y3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.250 0.805 1.51 1.26 ;
        RECT 1.250 0.805 2.875 0.87 ;
        RECT 2.620 0.090 2.88 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.115 0.630 0.83 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.055 0.090 1.705 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.915 0.090 2.37 0.74 ;
        END
    END c
END NAND3_Y3

MACRO NAND3_Y4
    CLASS CORE ;
    FOREIGN NAND3_Y4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.805 1.65 1.26 ;
        RECT 1.390 0.805 3.145 0.87 ;
        RECT 2.910 0.090 3.17 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.130 0.630 0.91 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.170 0.090 1.885 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.130 0.090 2.65 0.74 ;
        END
    END c
END NAND3_Y4

MACRO NAND3_Y6
    CLASS CORE ;
    FOREIGN NAND3_Y6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.805 1.995 1.26 ;
        RECT 1.670 0.805 3.815 0.87 ;
        RECT 3.490 0.090 3.815 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.155 0.630 1.065 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.405 0.090 2.25 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.555 0.090 3.14 0.74 ;
        END
    END c
END NAND3_Y6

MACRO NAND3_Y8
    CLASS CORE ;
    FOREIGN NAND3_Y8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.805 0.805 2.13 1.26 ;
        RECT 1.805 0.805 4.145 0.87 ;
        RECT 3.785 0.090 4.11 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.170 0.630 1.145 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.520 0.090 2.43 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.770 0.090 3.42 0.74 ;
        END
    END c
END NAND3_Y8

MACRO NAND3_Y10
    CLASS CORE ;
    FOREIGN NAND3_Y10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.805 2.475 1.26 ;
        RECT 2.085 0.805 4.75 0.87 ;
        RECT 4.365 0.090 4.755 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.195 0.630 1.365 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.755 0.090 2.795 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.195 0.090 3.975 0.74 ;
        END
    END c
END NAND3_Y10

MACRO NAND3_Y20
    CLASS CORE ;
    FOREIGN NAND3_Y20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.805 3.3 1.26 ;
        RECT 2.780 0.805 6.355 0.87 ;
        RECT 5.820 0.090 6.34 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.260 0.630 1.755 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.340 0.090 3.77 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.260 0.090 5.235 0.74 ;
        END
    END c
END NAND3_Y20

MACRO NAND3_Y40
    CLASS CORE ;
    FOREIGN NAND3_Y40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.890 0.805 4.605 1.26 ;
        RECT 3.890 0.805 8.895 0.87 ;
        RECT 8.150 0.090 8.865 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.365 0.630 2.51 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.275 0.090 5.225 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.965 0.090 7.395 0.74 ;
        END
    END c
END NAND3_Y40

MACRO NAND3_Y80
    CLASS CORE ;
    FOREIGN NAND3_Y80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.280 0.805 6.255 1.26 ;
        RECT 5.280 0.805 12.04 0.87 ;
        RECT 11.060 0.090 12.035 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.495 0.630 3.355 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.445 0.090 7.11 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.095 0.090 9.98 0.74 ;
        END
    END c
END NAND3_Y80

MACRO NAND3_Z1
    CLASS CORE ;
    FOREIGN NAND3_Z1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.415 0.805 0.48 1.26 ;
        RECT 0.415 0.805 0.935 0.87 ;
        RECT 0.875 0.090 0.94 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.040 0.630 0.3 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.350 0.090 0.545 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.640 0.090 0.77 0.74 ;
        END
    END c
END NAND3_Z1

MACRO NAND3_Z2
    CLASS CORE ;
    FOREIGN NAND3_Z2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.975 0.805 1.17 1.26 ;
        RECT 0.975 0.805 2.21 0.87 ;
        RECT 2.035 0.090 2.23 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.090 0.630 0.61 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.820 0.090 1.34 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.490 0.090 1.815 0.74 ;
        END
    END c
END NAND3_Z2

MACRO NAND3_Z3
    CLASS CORE ;
    FOREIGN NAND3_Z3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.250 0.805 1.51 1.26 ;
        RECT 1.250 0.805 2.875 0.87 ;
        RECT 2.620 0.090 2.88 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.115 0.630 0.83 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.055 0.090 1.705 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.915 0.090 2.37 0.74 ;
        END
    END c
END NAND3_Z3

MACRO NAND3_Z4
    CLASS CORE ;
    FOREIGN NAND3_Z4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.805 1.65 1.26 ;
        RECT 1.390 0.805 3.145 0.87 ;
        RECT 2.910 0.090 3.17 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.130 0.630 0.91 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.170 0.090 1.885 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.130 0.090 2.65 0.74 ;
        END
    END c
END NAND3_Z4

MACRO NAND3_Z6
    CLASS CORE ;
    FOREIGN NAND3_Z6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.805 1.995 1.26 ;
        RECT 1.670 0.805 3.815 0.87 ;
        RECT 3.490 0.090 3.815 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.155 0.630 1.065 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.405 0.090 2.25 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.555 0.090 3.14 0.74 ;
        END
    END c
END NAND3_Z6

MACRO NAND3_Z8
    CLASS CORE ;
    FOREIGN NAND3_Z8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.805 0.805 2.13 1.26 ;
        RECT 1.805 0.805 4.145 0.87 ;
        RECT 3.785 0.090 4.11 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.170 0.630 1.145 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.520 0.090 2.43 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.770 0.090 3.42 0.74 ;
        END
    END c
END NAND3_Z8

MACRO NAND3_Z10
    CLASS CORE ;
    FOREIGN NAND3_Z10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.805 2.475 1.26 ;
        RECT 2.085 0.805 4.75 0.87 ;
        RECT 4.365 0.090 4.755 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.195 0.630 1.365 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.755 0.090 2.795 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.195 0.090 3.975 0.74 ;
        END
    END c
END NAND3_Z10

MACRO NAND3_Z20
    CLASS CORE ;
    FOREIGN NAND3_Z20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.805 3.3 1.26 ;
        RECT 2.780 0.805 6.355 0.87 ;
        RECT 5.820 0.090 6.34 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.260 0.630 1.755 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.340 0.090 3.77 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.260 0.090 5.235 0.74 ;
        END
    END c
END NAND3_Z20

MACRO NAND3_Z40
    CLASS CORE ;
    FOREIGN NAND3_Z40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.890 0.805 4.605 1.26 ;
        RECT 3.890 0.805 8.895 0.87 ;
        RECT 8.150 0.090 8.865 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.365 0.630 2.51 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.275 0.090 5.225 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.965 0.090 7.395 0.74 ;
        END
    END c
END NAND3_Z40

MACRO NAND3_Z80
    CLASS CORE ;
    FOREIGN NAND3_Z80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.280 0.805 6.255 1.26 ;
        RECT 5.280 0.805 12.04 0.87 ;
        RECT 11.060 0.090 12.035 1.26 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.495 0.630 3.355 0.76 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.445 0.090 7.11 0.74 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.095 0.090 9.98 0.74 ;
        END
    END c
END NAND3_Z80

MACRO NAND4_X1
    CLASS CORE ;
    FOREIGN NAND4_X1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.210 0.53 0.925 ;
        RECT 0.465 0.870 0.79 0.935 ;
        RECT 0.715 0.870 0.78 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.725 1.34 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.725 1.085 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.635 0.405 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.725 0.83 0.79 ;
        END
    END d
END NAND4_X1

MACRO NAND4_X2
    CLASS CORE ;
    FOREIGN NAND4_X2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.040 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.210 1.12 0.925 ;
        RECT 0.925 0.870 1.575 0.935 ;
        RECT 1.435 0.870 1.63 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.285 0.725 2.61 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.780 0.725 2.105 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.635 0.745 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.725 1.6 0.79 ;
        END
    END d
END NAND4_X2

MACRO NAND4_X3
    CLASS CORE ;
    FOREIGN NAND4_X3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.210 1.355 0.925 ;
        RECT 1.160 0.870 2.005 0.935 ;
        RECT 1.790 0.870 1.985 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.860 0.725 3.25 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.225 0.725 2.615 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.635 0.915 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.590 0.725 1.98 0.79 ;
        END
    END d
END NAND4_X3

MACRO NAND4_X4
    CLASS CORE ;
    FOREIGN NAND4_X4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.210 1.65 0.925 ;
        RECT 1.390 0.870 2.43 0.935 ;
        RECT 2.150 0.870 2.41 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.430 0.725 3.95 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.725 3.19 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.635 1.15 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.910 0.725 2.43 0.79 ;
        END
    END d
END NAND4_X4

MACRO NAND4_X6
    CLASS CORE ;
    FOREIGN NAND4_X6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.210 1.945 0.925 ;
        RECT 1.620 0.870 2.79 0.935 ;
        RECT 2.510 0.870 2.835 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.725 4.585 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.725 3.7 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.635 1.32 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.725 2.815 0.79 ;
        END
    END d
END NAND4_X6

MACRO NAND4_X8
    CLASS CORE ;
    FOREIGN NAND4_X8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.210 2.18 0.925 ;
        RECT 1.855 0.870 3.22 0.935 ;
        RECT 2.865 0.870 3.19 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.725 5.225 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.725 4.21 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.840 0.635 1.49 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.725 3.195 0.79 ;
        END
    END d
END NAND4_X8

MACRO NAND4_X10
    CLASS CORE ;
    FOREIGN NAND4_X10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.970 0.210 2.36 0.925 ;
        RECT 1.970 0.870 3.4 0.935 ;
        RECT 3.045 0.870 3.435 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.860 0.725 5.575 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.785 0.725 4.5 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.895 0.635 1.61 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.705 0.725 3.42 0.79 ;
        END
    END d
END NAND4_X10

MACRO NAND4_X20
    CLASS CORE ;
    FOREIGN NAND4_X20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.665 0.210 3.185 0.925 ;
        RECT 2.665 0.870 4.615 0.935 ;
        RECT 4.120 0.870 4.64 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.575 0.725 7.55 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.115 0.725 6.09 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.210 0.635 2.185 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.660 0.725 4.635 0.79 ;
        END
    END d
END NAND4_X20

MACRO NAND4_X40
    CLASS CORE ;
    FOREIGN NAND4_X40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.210 4.24 0.925 ;
        RECT 3.590 0.870 6.255 0.935 ;
        RECT 5.555 0.870 6.205 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.860 0.725 10.16 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.895 0.725 8.195 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.625 0.635 2.925 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.935 0.725 6.235 0.79 ;
        END
    END d
END NAND4_X40

MACRO NAND4_X80
    CLASS CORE ;
    FOREIGN NAND4_X80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.340 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.980 0.210 5.89 0.925 ;
        RECT 4.980 0.870 8.62 0.935 ;
        RECT 7.705 0.870 8.615 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.290 0.725 14.11 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.565 0.725 11.385 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.255 0.635 4.075 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.845 0.725 8.665 0.79 ;
        END
    END d
END NAND4_X80

MACRO NAND4_Y1
    CLASS CORE ;
    FOREIGN NAND4_Y1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.210 0.53 0.925 ;
        RECT 0.465 0.870 0.79 0.935 ;
        RECT 0.715 0.870 0.78 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.725 1.34 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.725 1.085 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.635 0.405 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.725 0.83 0.79 ;
        END
    END d
END NAND4_Y1

MACRO NAND4_Y2
    CLASS CORE ;
    FOREIGN NAND4_Y2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.040 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.210 1.12 0.925 ;
        RECT 0.925 0.870 1.575 0.935 ;
        RECT 1.435 0.870 1.63 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.285 0.725 2.61 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.780 0.725 2.105 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.635 0.745 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.725 1.6 0.79 ;
        END
    END d
END NAND4_Y2

MACRO NAND4_Y3
    CLASS CORE ;
    FOREIGN NAND4_Y3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.210 1.355 0.925 ;
        RECT 1.160 0.870 2.005 0.935 ;
        RECT 1.790 0.870 1.985 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.860 0.725 3.25 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.225 0.725 2.615 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.635 0.915 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.590 0.725 1.98 0.79 ;
        END
    END d
END NAND4_Y3

MACRO NAND4_Y4
    CLASS CORE ;
    FOREIGN NAND4_Y4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.210 1.65 0.925 ;
        RECT 1.390 0.870 2.43 0.935 ;
        RECT 2.150 0.870 2.41 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.430 0.725 3.95 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.725 3.19 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.635 1.15 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.910 0.725 2.43 0.79 ;
        END
    END d
END NAND4_Y4

MACRO NAND4_Y6
    CLASS CORE ;
    FOREIGN NAND4_Y6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.210 1.945 0.925 ;
        RECT 1.620 0.870 2.79 0.935 ;
        RECT 2.510 0.870 2.835 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.725 4.585 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.725 3.7 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.635 1.32 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.725 2.815 0.79 ;
        END
    END d
END NAND4_Y6

MACRO NAND4_Y8
    CLASS CORE ;
    FOREIGN NAND4_Y8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.210 2.18 0.925 ;
        RECT 1.855 0.870 3.22 0.935 ;
        RECT 2.865 0.870 3.19 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.725 5.225 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.725 4.21 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.840 0.635 1.49 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.725 3.195 0.79 ;
        END
    END d
END NAND4_Y8

MACRO NAND4_Y10
    CLASS CORE ;
    FOREIGN NAND4_Y10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.970 0.210 2.36 0.925 ;
        RECT 1.970 0.870 3.4 0.935 ;
        RECT 3.045 0.870 3.435 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.860 0.725 5.575 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.785 0.725 4.5 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.895 0.635 1.61 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.705 0.725 3.42 0.79 ;
        END
    END d
END NAND4_Y10

MACRO NAND4_Y20
    CLASS CORE ;
    FOREIGN NAND4_Y20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.665 0.210 3.185 0.925 ;
        RECT 2.665 0.870 4.615 0.935 ;
        RECT 4.120 0.870 4.64 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.575 0.725 7.55 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.115 0.725 6.09 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.210 0.635 2.185 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.660 0.725 4.635 0.79 ;
        END
    END d
END NAND4_Y20

MACRO NAND4_Y40
    CLASS CORE ;
    FOREIGN NAND4_Y40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.210 4.24 0.925 ;
        RECT 3.590 0.870 6.255 0.935 ;
        RECT 5.555 0.870 6.205 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.860 0.725 10.16 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.895 0.725 8.195 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.625 0.635 2.925 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.935 0.725 6.235 0.79 ;
        END
    END d
END NAND4_Y40

MACRO NAND4_Y80
    CLASS CORE ;
    FOREIGN NAND4_Y80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.340 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.980 0.210 5.89 0.925 ;
        RECT 4.980 0.870 8.62 0.935 ;
        RECT 7.705 0.870 8.615 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.290 0.725 14.11 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.565 0.725 11.385 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.255 0.635 4.075 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.845 0.725 8.665 0.79 ;
        END
    END d
END NAND4_Y80

MACRO NAND4_Z1
    CLASS CORE ;
    FOREIGN NAND4_Z1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.210 0.53 0.925 ;
        RECT 0.465 0.870 0.79 0.935 ;
        RECT 0.715 0.870 0.78 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.725 1.34 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.725 1.085 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.210 0.635 0.405 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.725 0.83 0.79 ;
        END
    END d
END NAND4_Z1

MACRO NAND4_Z2
    CLASS CORE ;
    FOREIGN NAND4_Z2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.040 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.210 1.12 0.925 ;
        RECT 0.925 0.870 1.575 0.935 ;
        RECT 1.435 0.870 1.63 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.285 0.725 2.61 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.780 0.725 2.105 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.635 0.745 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.725 1.6 0.79 ;
        END
    END d
END NAND4_Z2

MACRO NAND4_Z3
    CLASS CORE ;
    FOREIGN NAND4_Z3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.210 1.355 0.925 ;
        RECT 1.160 0.870 2.005 0.935 ;
        RECT 1.790 0.870 1.985 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.860 0.725 3.25 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.225 0.725 2.615 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.525 0.635 0.915 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.590 0.725 1.98 0.79 ;
        END
    END d
END NAND4_Z3

MACRO NAND4_Z4
    CLASS CORE ;
    FOREIGN NAND4_Z4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.210 1.65 0.925 ;
        RECT 1.390 0.870 2.43 0.935 ;
        RECT 2.150 0.870 2.41 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.430 0.725 3.95 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.725 3.19 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.630 0.635 1.15 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.910 0.725 2.43 0.79 ;
        END
    END d
END NAND4_Z4

MACRO NAND4_Z6
    CLASS CORE ;
    FOREIGN NAND4_Z6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.210 1.945 0.925 ;
        RECT 1.620 0.870 2.79 0.935 ;
        RECT 2.510 0.870 2.835 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.725 4.585 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.725 3.7 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.735 0.635 1.32 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.725 2.815 0.79 ;
        END
    END d
END NAND4_Z6

MACRO NAND4_Z8
    CLASS CORE ;
    FOREIGN NAND4_Z8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.210 2.18 0.925 ;
        RECT 1.855 0.870 3.22 0.935 ;
        RECT 2.865 0.870 3.19 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.725 5.225 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.725 4.21 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.840 0.635 1.49 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.725 3.195 0.79 ;
        END
    END d
END NAND4_Z8

MACRO NAND4_Z10
    CLASS CORE ;
    FOREIGN NAND4_Z10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.970 0.210 2.36 0.925 ;
        RECT 1.970 0.870 3.4 0.935 ;
        RECT 3.045 0.870 3.435 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.860 0.725 5.575 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.785 0.725 4.5 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.895 0.635 1.61 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.705 0.725 3.42 0.79 ;
        END
    END d
END NAND4_Z10

MACRO NAND4_Z20
    CLASS CORE ;
    FOREIGN NAND4_Z20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.665 0.210 3.185 0.925 ;
        RECT 2.665 0.870 4.615 0.935 ;
        RECT 4.120 0.870 4.64 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.575 0.725 7.55 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.115 0.725 6.09 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.210 0.635 2.185 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.660 0.725 4.635 0.79 ;
        END
    END d
END NAND4_Z20

MACRO NAND4_Z40
    CLASS CORE ;
    FOREIGN NAND4_Z40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.210 4.24 0.925 ;
        RECT 3.590 0.870 6.255 0.935 ;
        RECT 5.555 0.870 6.205 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.860 0.725 10.16 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.895 0.725 8.195 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.625 0.635 2.925 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.935 0.725 6.235 0.79 ;
        END
    END d
END NAND4_Z40

MACRO NAND4_Z80
    CLASS CORE ;
    FOREIGN NAND4_Z80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.340 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.980 0.210 5.89 0.925 ;
        RECT 4.980 0.870 8.62 0.935 ;
        RECT 7.705 0.870 8.615 1.52 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.290 0.725 14.11 0.79 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.565 0.725 11.385 0.79 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.255 0.635 4.075 0.7 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.845 0.725 8.665 0.79 ;
        END
    END d
END NAND4_Z80

MACRO NOR2_X1
    CLASS CORE ;
    FOREIGN NOR2_X1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.520 0.150 0.65 0.54 ;
        RECT 0.465 0.150 0.66 0.28 ;
        RECT 0.520 0.505 0.91 0.57 ;
        RECT 0.805 0.505 0.935 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.235 0.340 0.43 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.715 0.340 0.91 0.405 ;
        END
    END b
END NOR2_X1

MACRO NOR2_X2
    CLASS CORE ;
    FOREIGN NOR2_X2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.215 0.150 1.475 0.54 ;
        RECT 1.085 0.150 1.54 0.28 ;
        RECT 1.215 0.505 2.125 0.57 ;
        RECT 1.875 0.505 2.135 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.550 0.340 1.005 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.340 2.125 0.405 ;
        END
    END b
END NOR2_X2

MACRO NOR2_X3
    CLASS CORE ;
    FOREIGN NOR2_X3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.565 0.150 1.89 0.54 ;
        RECT 1.395 0.150 1.98 0.28 ;
        RECT 1.565 0.505 2.67 0.57 ;
        RECT 2.410 0.505 2.735 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.710 0.340 1.295 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.340 2.735 0.405 ;
        END
    END b
END NOR2_X3

MACRO NOR2_X4
    CLASS CORE ;
    FOREIGN NOR2_X4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.740 0.150 2.065 0.54 ;
        RECT 1.550 0.150 2.2 0.28 ;
        RECT 1.740 0.505 2.975 0.57 ;
        RECT 2.675 0.505 3.0 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.790 0.340 1.44 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.390 0.340 3.04 0.405 ;
        END
    END b
END NOR2_X4

MACRO NOR2_X6
    CLASS CORE ;
    FOREIGN NOR2_X6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.150 2.475 0.54 ;
        RECT 1.860 0.150 2.64 0.28 ;
        RECT 2.085 0.505 3.58 0.57 ;
        RECT 3.210 0.505 3.6 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.945 0.340 1.725 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.865 0.340 3.645 0.405 ;
        END
    END b
END NOR2_X6

MACRO NOR2_X8
    CLASS CORE ;
    FOREIGN NOR2_X8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.260 0.150 2.715 0.54 ;
        RECT 2.015 0.150 2.86 0.28 ;
        RECT 2.260 0.505 3.885 0.57 ;
        RECT 3.480 0.505 3.935 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.025 0.340 1.87 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.105 0.340 3.95 0.405 ;
        END
    END b
END NOR2_X8

MACRO NOR2_X10
    CLASS CORE ;
    FOREIGN NOR2_X10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.605 0.150 3.125 0.54 ;
        RECT 2.325 0.150 3.365 0.28 ;
        RECT 2.605 0.505 4.49 0.57 ;
        RECT 4.015 0.505 4.535 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.180 0.340 2.09 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.580 0.340 4.49 0.405 ;
        END
    END b
END NOR2_X10

MACRO NOR2_X20
    CLASS CORE ;
    FOREIGN NOR2_X20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.475 0.150 4.125 0.54 ;
        RECT 3.100 0.150 4.465 0.28 ;
        RECT 3.475 0.505 6.01 0.57 ;
        RECT 5.350 0.505 6.0 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.575 0.340 2.81 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.775 0.340 6.01 0.405 ;
        END
    END b
END NOR2_X20

MACRO NOR2_X40
    CLASS CORE ;
    FOREIGN NOR2_X40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.865 0.150 5.775 0.54 ;
        RECT 4.340 0.150 6.225 0.28 ;
        RECT 4.865 0.505 8.375 0.57 ;
        RECT 7.490 0.505 8.4 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.205 0.340 3.96 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.685 0.340 8.44 0.405 ;
        END
    END b
END NOR2_X40

MACRO NOR2_X80
    CLASS CORE ;
    FOREIGN NOR2_X80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.605 0.150 7.84 0.54 ;
        RECT 5.890 0.150 8.425 0.28 ;
        RECT 6.605 0.505 11.415 0.57 ;
        RECT 10.165 0.505 11.4 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.995 0.340 5.4 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.075 0.340 11.48 0.405 ;
        END
    END b
END NOR2_X80

MACRO NOR2_Y1
    CLASS CORE ;
    FOREIGN NOR2_Y1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.520 0.150 0.65 0.54 ;
        RECT 0.465 0.150 0.66 0.28 ;
        RECT 0.520 0.505 0.91 0.57 ;
        RECT 0.805 0.505 0.935 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.235 0.340 0.43 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.715 0.340 0.91 0.405 ;
        END
    END b
END NOR2_Y1

MACRO NOR2_Y2
    CLASS CORE ;
    FOREIGN NOR2_Y2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.215 0.150 1.475 0.54 ;
        RECT 1.085 0.150 1.54 0.28 ;
        RECT 1.215 0.505 2.125 0.57 ;
        RECT 1.875 0.505 2.135 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.550 0.340 1.005 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.340 2.125 0.405 ;
        END
    END b
END NOR2_Y2

MACRO NOR2_Y3
    CLASS CORE ;
    FOREIGN NOR2_Y3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.565 0.150 1.89 0.54 ;
        RECT 1.395 0.150 1.98 0.28 ;
        RECT 1.565 0.505 2.67 0.57 ;
        RECT 2.410 0.505 2.735 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.710 0.340 1.295 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.340 2.735 0.405 ;
        END
    END b
END NOR2_Y3

MACRO NOR2_Y4
    CLASS CORE ;
    FOREIGN NOR2_Y4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.740 0.150 2.065 0.54 ;
        RECT 1.550 0.150 2.2 0.28 ;
        RECT 1.740 0.505 2.975 0.57 ;
        RECT 2.675 0.505 3.0 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.790 0.340 1.44 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.390 0.340 3.04 0.405 ;
        END
    END b
END NOR2_Y4

MACRO NOR2_Y6
    CLASS CORE ;
    FOREIGN NOR2_Y6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.150 2.475 0.54 ;
        RECT 1.860 0.150 2.64 0.28 ;
        RECT 2.085 0.505 3.58 0.57 ;
        RECT 3.210 0.505 3.6 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.945 0.340 1.725 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.865 0.340 3.645 0.405 ;
        END
    END b
END NOR2_Y6

MACRO NOR2_Y8
    CLASS CORE ;
    FOREIGN NOR2_Y8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.260 0.150 2.715 0.54 ;
        RECT 2.015 0.150 2.86 0.28 ;
        RECT 2.260 0.505 3.885 0.57 ;
        RECT 3.480 0.505 3.935 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.025 0.340 1.87 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.105 0.340 3.95 0.405 ;
        END
    END b
END NOR2_Y8

MACRO NOR2_Y10
    CLASS CORE ;
    FOREIGN NOR2_Y10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.605 0.150 3.125 0.54 ;
        RECT 2.325 0.150 3.365 0.28 ;
        RECT 2.605 0.505 4.49 0.57 ;
        RECT 4.015 0.505 4.535 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.180 0.340 2.09 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.580 0.340 4.49 0.405 ;
        END
    END b
END NOR2_Y10

MACRO NOR2_Y20
    CLASS CORE ;
    FOREIGN NOR2_Y20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.475 0.150 4.125 0.54 ;
        RECT 3.100 0.150 4.465 0.28 ;
        RECT 3.475 0.505 6.01 0.57 ;
        RECT 5.350 0.505 6.0 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.575 0.340 2.81 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.775 0.340 6.01 0.405 ;
        END
    END b
END NOR2_Y20

MACRO NOR2_Y40
    CLASS CORE ;
    FOREIGN NOR2_Y40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.865 0.150 5.775 0.54 ;
        RECT 4.340 0.150 6.225 0.28 ;
        RECT 4.865 0.505 8.375 0.57 ;
        RECT 7.490 0.505 8.4 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.205 0.340 3.96 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.685 0.340 8.44 0.405 ;
        END
    END b
END NOR2_Y40

MACRO NOR2_Y80
    CLASS CORE ;
    FOREIGN NOR2_Y80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.605 0.150 7.84 0.54 ;
        RECT 5.890 0.150 8.425 0.28 ;
        RECT 6.605 0.505 11.415 0.57 ;
        RECT 10.165 0.505 11.4 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.995 0.340 5.4 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.075 0.340 11.48 0.405 ;
        END
    END b
END NOR2_Y80

MACRO NOR2_Z1
    CLASS CORE ;
    FOREIGN NOR2_Z1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.520 0.150 0.65 0.54 ;
        RECT 0.465 0.150 0.66 0.28 ;
        RECT 0.520 0.505 0.91 0.57 ;
        RECT 0.805 0.505 0.935 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.235 0.340 0.43 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.715 0.340 0.91 0.405 ;
        END
    END b
END NOR2_Z1

MACRO NOR2_Z2
    CLASS CORE ;
    FOREIGN NOR2_Z2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.215 0.150 1.475 0.54 ;
        RECT 1.085 0.150 1.54 0.28 ;
        RECT 1.215 0.505 2.125 0.57 ;
        RECT 1.875 0.505 2.135 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.550 0.340 1.005 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.340 2.125 0.405 ;
        END
    END b
END NOR2_Z2

MACRO NOR2_Z3
    CLASS CORE ;
    FOREIGN NOR2_Z3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.565 0.150 1.89 0.54 ;
        RECT 1.395 0.150 1.98 0.28 ;
        RECT 1.565 0.505 2.67 0.57 ;
        RECT 2.410 0.505 2.735 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.710 0.340 1.295 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.340 2.735 0.405 ;
        END
    END b
END NOR2_Z3

MACRO NOR2_Z4
    CLASS CORE ;
    FOREIGN NOR2_Z4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.740 0.150 2.065 0.54 ;
        RECT 1.550 0.150 2.2 0.28 ;
        RECT 1.740 0.505 2.975 0.57 ;
        RECT 2.675 0.505 3.0 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.790 0.340 1.44 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.390 0.340 3.04 0.405 ;
        END
    END b
END NOR2_Z4

MACRO NOR2_Z6
    CLASS CORE ;
    FOREIGN NOR2_Z6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.150 2.475 0.54 ;
        RECT 1.860 0.150 2.64 0.28 ;
        RECT 2.085 0.505 3.58 0.57 ;
        RECT 3.210 0.505 3.6 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.945 0.340 1.725 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.865 0.340 3.645 0.405 ;
        END
    END b
END NOR2_Z6

MACRO NOR2_Z8
    CLASS CORE ;
    FOREIGN NOR2_Z8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.260 0.150 2.715 0.54 ;
        RECT 2.015 0.150 2.86 0.28 ;
        RECT 2.260 0.505 3.885 0.57 ;
        RECT 3.480 0.505 3.935 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.025 0.340 1.87 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.105 0.340 3.95 0.405 ;
        END
    END b
END NOR2_Z8

MACRO NOR2_Z10
    CLASS CORE ;
    FOREIGN NOR2_Z10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.605 0.150 3.125 0.54 ;
        RECT 2.325 0.150 3.365 0.28 ;
        RECT 2.605 0.505 4.49 0.57 ;
        RECT 4.015 0.505 4.535 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.180 0.340 2.09 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.580 0.340 4.49 0.405 ;
        END
    END b
END NOR2_Z10

MACRO NOR2_Z20
    CLASS CORE ;
    FOREIGN NOR2_Z20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.475 0.150 4.125 0.54 ;
        RECT 3.100 0.150 4.465 0.28 ;
        RECT 3.475 0.505 6.01 0.57 ;
        RECT 5.350 0.505 6.0 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.575 0.340 2.81 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.775 0.340 6.01 0.405 ;
        END
    END b
END NOR2_Z20

MACRO NOR2_Z40
    CLASS CORE ;
    FOREIGN NOR2_Z40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.865 0.150 5.775 0.54 ;
        RECT 4.340 0.150 6.225 0.28 ;
        RECT 4.865 0.505 8.375 0.57 ;
        RECT 7.490 0.505 8.4 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.205 0.340 3.96 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.685 0.340 8.44 0.405 ;
        END
    END b
END NOR2_Z40

MACRO NOR2_Z80
    CLASS CORE ;
    FOREIGN NOR2_Z80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.605 0.150 7.84 0.54 ;
        RECT 5.890 0.150 8.425 0.28 ;
        RECT 6.605 0.505 11.415 0.57 ;
        RECT 10.165 0.505 11.4 1.155 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.995 0.340 5.4 0.405 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.075 0.340 11.48 0.405 ;
        END
    END b
END NOR2_Z80

MACRO NOR3_X1
    CLASS CORE ;
    FOREIGN NOR3_X1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.130 0.485 0.39 ;
        RECT 0.420 0.340 0.94 0.405 ;
        RECT 0.870 0.130 0.935 1.625 ;
        RECT 0.870 0.545 0.935 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.085 0.365 0.28 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.415 0.430 0.545 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.645 0.430 0.775 0.56 ;
        END
    END c
END NOR3_X1

MACRO NOR3_X2
    CLASS CORE ;
    FOREIGN NOR3_X2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.980 0.130 1.175 0.39 ;
        RECT 0.980 0.340 2.215 0.405 ;
        RECT 2.030 0.130 2.225 1.625 ;
        RECT 2.030 0.545 2.225 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.195 0.365 0.65 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.975 0.430 1.3 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.505 0.430 1.83 0.56 ;
        END
    END c
END NOR3_X2

MACRO NOR3_X3
    CLASS CORE ;
    FOREIGN NOR3_X3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.260 0.130 1.52 0.39 ;
        RECT 1.260 0.340 2.82 0.405 ;
        RECT 2.610 0.130 2.87 1.625 ;
        RECT 2.610 0.545 2.87 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.365 0.77 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.250 0.430 1.705 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.935 0.430 2.39 0.56 ;
        END
    END c
END NOR3_X3

MACRO NOR3_X4
    CLASS CORE ;
    FOREIGN NOR3_X4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.400 0.130 1.66 0.39 ;
        RECT 1.400 0.340 3.155 0.405 ;
        RECT 2.900 0.130 3.16 1.625 ;
        RECT 2.900 0.545 3.16 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.280 0.365 0.865 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.430 1.845 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.430 2.67 0.56 ;
        END
    END c
END NOR3_X4

MACRO NOR3_X6
    CLASS CORE ;
    FOREIGN NOR3_X6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.680 0.130 2.005 0.39 ;
        RECT 1.680 0.340 3.76 0.405 ;
        RECT 3.480 0.130 3.805 1.625 ;
        RECT 3.480 0.545 3.805 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.335 0.365 1.05 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.430 2.255 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.430 3.165 0.56 ;
        END
    END c
END NOR3_X6

MACRO NOR3_X8
    CLASS CORE ;
    FOREIGN NOR3_X8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.820 0.130 2.145 0.39 ;
        RECT 1.820 0.340 4.095 0.405 ;
        RECT 3.770 0.130 4.095 1.625 ;
        RECT 3.770 0.545 4.095 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.365 0.365 1.145 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.805 0.430 2.39 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.795 0.430 3.445 0.56 ;
        END
    END c
END NOR3_X8

MACRO NOR3_X10
    CLASS CORE ;
    FOREIGN NOR3_X10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.100 0.130 2.49 0.39 ;
        RECT 2.100 0.340 4.765 0.405 ;
        RECT 4.350 0.130 4.74 1.625 ;
        RECT 4.350 0.545 4.74 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.365 1.33 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.430 2.8 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.225 0.430 3.94 0.56 ;
        END
    END c
END NOR3_X10

MACRO NOR3_X20
    CLASS CORE ;
    FOREIGN NOR3_X20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.800 0.130 3.32 0.39 ;
        RECT 2.800 0.340 6.31 0.405 ;
        RECT 5.800 0.130 6.32 1.625 ;
        RECT 5.800 0.545 6.32 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.560 0.365 1.795 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.430 3.69 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.430 5.275 0.56 ;
        END
    END c
END NOR3_X20

MACRO NOR3_X40
    CLASS CORE ;
    FOREIGN NOR3_X40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.920 0.130 4.635 0.39 ;
        RECT 3.920 0.340 8.86 0.405 ;
        RECT 8.120 0.130 8.835 1.625 ;
        RECT 8.120 0.545 8.9 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.785 0.365 2.475 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.890 0.430 5.19 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.020 0.430 7.385 0.56 ;
        END
    END c
END NOR3_X40

MACRO NOR3_X80
    CLASS CORE ;
    FOREIGN NOR3_X80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.320 0.130 6.295 0.39 ;
        RECT 5.320 0.340 12.015 0.405 ;
        RECT 11.020 0.130 11.995 1.625 ;
        RECT 11.020 0.545 12.06 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.065 0.365 3.405 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.280 0.430 7.035 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.170 0.430 10.055 0.56 ;
        END
    END c
END NOR3_X80

MACRO NOR3_Y1
    CLASS CORE ;
    FOREIGN NOR3_Y1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.130 0.485 0.39 ;
        RECT 0.420 0.340 0.94 0.405 ;
        RECT 0.870 0.130 0.935 1.625 ;
        RECT 0.870 0.545 0.935 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.085 0.365 0.28 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.415 0.430 0.545 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.645 0.430 0.775 0.56 ;
        END
    END c
END NOR3_Y1

MACRO NOR3_Y2
    CLASS CORE ;
    FOREIGN NOR3_Y2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.980 0.130 1.175 0.39 ;
        RECT 0.980 0.340 2.215 0.405 ;
        RECT 2.030 0.130 2.225 1.625 ;
        RECT 2.030 0.545 2.225 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.195 0.365 0.65 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.975 0.430 1.3 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.505 0.430 1.83 0.56 ;
        END
    END c
END NOR3_Y2

MACRO NOR3_Y3
    CLASS CORE ;
    FOREIGN NOR3_Y3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.260 0.130 1.52 0.39 ;
        RECT 1.260 0.340 2.82 0.405 ;
        RECT 2.610 0.130 2.87 1.625 ;
        RECT 2.610 0.545 2.87 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.365 0.77 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.250 0.430 1.705 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.935 0.430 2.39 0.56 ;
        END
    END c
END NOR3_Y3

MACRO NOR3_Y4
    CLASS CORE ;
    FOREIGN NOR3_Y4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.400 0.130 1.66 0.39 ;
        RECT 1.400 0.340 3.155 0.405 ;
        RECT 2.900 0.130 3.16 1.625 ;
        RECT 2.900 0.545 3.16 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.280 0.365 0.865 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.430 1.845 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.430 2.67 0.56 ;
        END
    END c
END NOR3_Y4

MACRO NOR3_Y6
    CLASS CORE ;
    FOREIGN NOR3_Y6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.680 0.130 2.005 0.39 ;
        RECT 1.680 0.340 3.76 0.405 ;
        RECT 3.480 0.130 3.805 1.625 ;
        RECT 3.480 0.545 3.805 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.335 0.365 1.05 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.430 2.255 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.430 3.165 0.56 ;
        END
    END c
END NOR3_Y6

MACRO NOR3_Y8
    CLASS CORE ;
    FOREIGN NOR3_Y8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.820 0.130 2.145 0.39 ;
        RECT 1.820 0.340 4.095 0.405 ;
        RECT 3.770 0.130 4.095 1.625 ;
        RECT 3.770 0.545 4.095 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.365 0.365 1.145 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.805 0.430 2.39 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.795 0.430 3.445 0.56 ;
        END
    END c
END NOR3_Y8

MACRO NOR3_Y10
    CLASS CORE ;
    FOREIGN NOR3_Y10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.100 0.130 2.49 0.39 ;
        RECT 2.100 0.340 4.765 0.405 ;
        RECT 4.350 0.130 4.74 1.625 ;
        RECT 4.350 0.545 4.74 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.365 1.33 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.430 2.8 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.225 0.430 3.94 0.56 ;
        END
    END c
END NOR3_Y10

MACRO NOR3_Y20
    CLASS CORE ;
    FOREIGN NOR3_Y20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.800 0.130 3.32 0.39 ;
        RECT 2.800 0.340 6.31 0.405 ;
        RECT 5.800 0.130 6.32 1.625 ;
        RECT 5.800 0.545 6.32 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.560 0.365 1.795 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.430 3.69 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.430 5.275 0.56 ;
        END
    END c
END NOR3_Y20

MACRO NOR3_Y40
    CLASS CORE ;
    FOREIGN NOR3_Y40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.920 0.130 4.635 0.39 ;
        RECT 3.920 0.340 8.86 0.405 ;
        RECT 8.120 0.130 8.835 1.625 ;
        RECT 8.120 0.545 8.9 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.785 0.365 2.475 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.890 0.430 5.19 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.020 0.430 7.385 0.56 ;
        END
    END c
END NOR3_Y40

MACRO NOR3_Y80
    CLASS CORE ;
    FOREIGN NOR3_Y80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.320 0.130 6.295 0.39 ;
        RECT 5.320 0.340 12.015 0.405 ;
        RECT 11.020 0.130 11.995 1.625 ;
        RECT 11.020 0.545 12.06 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.065 0.365 3.405 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.280 0.430 7.035 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.170 0.430 10.055 0.56 ;
        END
    END c
END NOR3_Y80

MACRO NOR3_Z1
    CLASS CORE ;
    FOREIGN NOR3_Z1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.140 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.130 0.485 0.39 ;
        RECT 0.420 0.340 0.94 0.405 ;
        RECT 0.870 0.130 0.935 1.625 ;
        RECT 0.870 0.545 0.935 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.085 0.365 0.28 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.415 0.430 0.545 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.645 0.430 0.775 0.56 ;
        END
    END c
END NOR3_Z1

MACRO NOR3_Z2
    CLASS CORE ;
    FOREIGN NOR3_Z2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 2.660 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.980 0.130 1.175 0.39 ;
        RECT 0.980 0.340 2.215 0.405 ;
        RECT 2.030 0.130 2.225 1.625 ;
        RECT 2.030 0.545 2.225 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.195 0.365 0.65 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.975 0.430 1.3 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.505 0.430 1.83 0.56 ;
        END
    END c
END NOR3_Z2

MACRO NOR3_Z3
    CLASS CORE ;
    FOREIGN NOR3_Z3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.420 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.260 0.130 1.52 0.39 ;
        RECT 1.260 0.340 2.82 0.405 ;
        RECT 2.610 0.130 2.87 1.625 ;
        RECT 2.610 0.545 2.87 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.365 0.77 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.250 0.430 1.705 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.935 0.430 2.39 0.56 ;
        END
    END c
END NOR3_Z3

MACRO NOR3_Z4
    CLASS CORE ;
    FOREIGN NOR3_Z4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.400 0.130 1.66 0.39 ;
        RECT 1.400 0.340 3.155 0.405 ;
        RECT 2.900 0.130 3.16 1.625 ;
        RECT 2.900 0.545 3.16 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.280 0.365 0.865 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.430 1.845 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.150 0.430 2.67 0.56 ;
        END
    END c
END NOR3_Z4

MACRO NOR3_Z6
    CLASS CORE ;
    FOREIGN NOR3_Z6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.680 0.130 2.005 0.39 ;
        RECT 1.680 0.340 3.76 0.405 ;
        RECT 3.480 0.130 3.805 1.625 ;
        RECT 3.480 0.545 3.805 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.335 0.365 1.05 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.670 0.430 2.255 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.580 0.430 3.165 0.56 ;
        END
    END c
END NOR3_Z6

MACRO NOR3_Z8
    CLASS CORE ;
    FOREIGN NOR3_Z8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.940 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.820 0.130 2.145 0.39 ;
        RECT 1.820 0.340 4.095 0.405 ;
        RECT 3.770 0.130 4.095 1.625 ;
        RECT 3.770 0.545 4.095 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.365 0.365 1.145 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.805 0.430 2.39 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.795 0.430 3.445 0.56 ;
        END
    END c
END NOR3_Z8

MACRO NOR3_Z10
    CLASS CORE ;
    FOREIGN NOR3_Z10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.700 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.100 0.130 2.49 0.39 ;
        RECT 2.100 0.340 4.765 0.405 ;
        RECT 4.350 0.130 4.74 1.625 ;
        RECT 4.350 0.545 4.74 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.420 0.365 1.33 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.085 0.430 2.8 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.225 0.430 3.94 0.56 ;
        END
    END c
END NOR3_Z10

MACRO NOR3_Z20
    CLASS CORE ;
    FOREIGN NOR3_Z20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 7.600 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.800 0.130 3.32 0.39 ;
        RECT 2.800 0.340 6.31 0.405 ;
        RECT 5.800 0.130 6.32 1.625 ;
        RECT 5.800 0.545 6.32 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.560 0.365 1.795 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.780 0.430 3.69 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.300 0.430 5.275 0.56 ;
        END
    END c
END NOR3_Z20

MACRO NOR3_Z40
    CLASS CORE ;
    FOREIGN NOR3_Z40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 10.640 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.920 0.130 4.635 0.39 ;
        RECT 3.920 0.340 8.86 0.405 ;
        RECT 8.120 0.130 8.835 1.625 ;
        RECT 8.120 0.545 8.9 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.785 0.365 2.475 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.890 0.430 5.19 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.020 0.430 7.385 0.56 ;
        END
    END c
END NOR3_Z40

MACRO NOR3_Z80
    CLASS CORE ;
    FOREIGN NOR3_Z80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 14.440 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.320 0.130 6.295 0.39 ;
        RECT 5.320 0.340 12.015 0.405 ;
        RECT 11.020 0.130 11.995 1.625 ;
        RECT 11.020 0.545 12.06 1.585 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.065 0.365 3.405 0.43 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.280 0.430 7.035 0.56 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.170 0.430 10.055 0.56 ;
        END
    END c
END NOR3_Z80

MACRO NOR4_X1
    CLASS CORE ;
    FOREIGN NOR4_X1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.090 0.53 1.455 ;
        RECT 0.465 0.090 0.79 0.155 ;
        RECT 0.715 0.090 0.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.530 1.34 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.530 1.085 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.045 0.530 0.305 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.530 0.83 0.66 ;
        END
    END d
END NOR4_X1

MACRO NOR4_X2
    CLASS CORE ;
    FOREIGN NOR4_X2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.040 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.090 1.12 1.455 ;
        RECT 0.925 0.090 1.575 0.155 ;
        RECT 1.425 0.090 1.62 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.285 0.530 2.61 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.780 0.530 2.105 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.085 0.530 0.605 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.530 1.6 0.66 ;
        END
    END d
END NOR4_X2

MACRO NOR4_X3
    CLASS CORE ;
    FOREIGN NOR4_X3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.090 1.355 1.455 ;
        RECT 1.160 0.090 2.005 0.155 ;
        RECT 1.785 0.090 1.98 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.860 0.530 3.25 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.225 0.530 2.615 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.110 0.530 0.76 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.590 0.530 1.98 0.66 ;
        END
    END d
END NOR4_X3

MACRO NOR4_X4
    CLASS CORE ;
    FOREIGN NOR4_X4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.090 1.65 1.455 ;
        RECT 1.390 0.090 2.43 0.155 ;
        RECT 2.140 0.090 2.4 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.430 0.530 3.95 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.530 3.19 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.130 0.530 0.91 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.910 0.530 2.43 0.66 ;
        END
    END d
END NOR4_X4

MACRO NOR4_X6
    CLASS CORE ;
    FOREIGN NOR4_X6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.090 1.945 1.455 ;
        RECT 1.620 0.090 2.79 0.155 ;
        RECT 2.495 0.090 2.82 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.530 4.585 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.530 3.7 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.150 0.530 1.06 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.530 2.815 0.66 ;
        END
    END d
END NOR4_X6

MACRO NOR4_X8
    CLASS CORE ;
    FOREIGN NOR4_X8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.090 2.18 1.455 ;
        RECT 1.855 0.090 3.22 0.155 ;
        RECT 2.855 0.090 3.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.530 5.225 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.530 4.21 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.175 0.530 1.215 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.530 3.195 0.66 ;
        END
    END d
END NOR4_X8

MACRO NOR4_X10
    CLASS CORE ;
    FOREIGN NOR4_X10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.970 0.090 2.36 1.455 ;
        RECT 1.970 0.090 3.4 0.155 ;
        RECT 3.030 0.090 3.42 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.860 0.530 5.575 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.785 0.530 4.5 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.185 0.530 1.29 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.705 0.530 3.42 0.66 ;
        END
    END d
END NOR4_X10

MACRO NOR4_X20
    CLASS CORE ;
    FOREIGN NOR4_X20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.665 0.090 3.185 1.455 ;
        RECT 2.665 0.090 4.615 0.155 ;
        RECT 4.100 0.090 4.62 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.575 0.530 7.55 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.115 0.530 6.09 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.530 1.68 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.660 0.530 4.635 0.66 ;
        END
    END d
END NOR4_X20

MACRO NOR4_X40
    CLASS CORE ;
    FOREIGN NOR4_X40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.090 4.24 1.455 ;
        RECT 3.590 0.090 6.19 0.155 ;
        RECT 5.530 0.090 6.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.860 0.530 10.16 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.895 0.530 8.195 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.335 0.530 2.285 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.935 0.530 6.235 0.66 ;
        END
    END d
END NOR4_X40

MACRO NOR4_X80
    CLASS CORE ;
    FOREIGN NOR4_X80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.340 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.980 0.090 5.89 1.455 ;
        RECT 4.980 0.090 8.62 0.155 ;
        RECT 7.670 0.090 8.58 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.290 0.530 14.11 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.565 0.530 11.385 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.530 3.195 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.845 0.530 8.665 0.66 ;
        END
    END d
END NOR4_X80

MACRO NOR4_Y1
    CLASS CORE ;
    FOREIGN NOR4_Y1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.090 0.53 1.455 ;
        RECT 0.465 0.090 0.79 0.155 ;
        RECT 0.715 0.090 0.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.530 1.34 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.530 1.085 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.045 0.530 0.305 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.530 0.83 0.66 ;
        END
    END d
END NOR4_Y1

MACRO NOR4_Y2
    CLASS CORE ;
    FOREIGN NOR4_Y2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.040 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.090 1.12 1.455 ;
        RECT 0.925 0.090 1.575 0.155 ;
        RECT 1.425 0.090 1.62 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.285 0.530 2.61 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.780 0.530 2.105 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.085 0.530 0.605 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.530 1.6 0.66 ;
        END
    END d
END NOR4_Y2

MACRO NOR4_Y3
    CLASS CORE ;
    FOREIGN NOR4_Y3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.090 1.355 1.455 ;
        RECT 1.160 0.090 2.005 0.155 ;
        RECT 1.785 0.090 1.98 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.860 0.530 3.25 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.225 0.530 2.615 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.110 0.530 0.76 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.590 0.530 1.98 0.66 ;
        END
    END d
END NOR4_Y3

MACRO NOR4_Y4
    CLASS CORE ;
    FOREIGN NOR4_Y4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.090 1.65 1.455 ;
        RECT 1.390 0.090 2.43 0.155 ;
        RECT 2.140 0.090 2.4 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.430 0.530 3.95 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.530 3.19 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.130 0.530 0.91 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.910 0.530 2.43 0.66 ;
        END
    END d
END NOR4_Y4

MACRO NOR4_Y6
    CLASS CORE ;
    FOREIGN NOR4_Y6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.090 1.945 1.455 ;
        RECT 1.620 0.090 2.79 0.155 ;
        RECT 2.495 0.090 2.82 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.530 4.585 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.530 3.7 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.150 0.530 1.06 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.530 2.815 0.66 ;
        END
    END d
END NOR4_Y6

MACRO NOR4_Y8
    CLASS CORE ;
    FOREIGN NOR4_Y8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.090 2.18 1.455 ;
        RECT 1.855 0.090 3.22 0.155 ;
        RECT 2.855 0.090 3.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.530 5.225 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.530 4.21 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.175 0.530 1.215 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.530 3.195 0.66 ;
        END
    END d
END NOR4_Y8

MACRO NOR4_Y10
    CLASS CORE ;
    FOREIGN NOR4_Y10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.970 0.090 2.36 1.455 ;
        RECT 1.970 0.090 3.4 0.155 ;
        RECT 3.030 0.090 3.42 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.860 0.530 5.575 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.785 0.530 4.5 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.185 0.530 1.29 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.705 0.530 3.42 0.66 ;
        END
    END d
END NOR4_Y10

MACRO NOR4_Y20
    CLASS CORE ;
    FOREIGN NOR4_Y20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.665 0.090 3.185 1.455 ;
        RECT 2.665 0.090 4.615 0.155 ;
        RECT 4.100 0.090 4.62 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.575 0.530 7.55 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.115 0.530 6.09 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.530 1.68 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.660 0.530 4.635 0.66 ;
        END
    END d
END NOR4_Y20

MACRO NOR4_Y40
    CLASS CORE ;
    FOREIGN NOR4_Y40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.090 4.24 1.455 ;
        RECT 3.590 0.090 6.19 0.155 ;
        RECT 5.530 0.090 6.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.860 0.530 10.16 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.895 0.530 8.195 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.335 0.530 2.285 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.935 0.530 6.235 0.66 ;
        END
    END d
END NOR4_Y40

MACRO NOR4_Y80
    CLASS CORE ;
    FOREIGN NOR4_Y80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.340 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.980 0.090 5.89 1.455 ;
        RECT 4.980 0.090 8.62 0.155 ;
        RECT 7.670 0.090 8.58 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.290 0.530 14.11 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.565 0.530 11.385 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.530 3.195 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.845 0.530 8.665 0.66 ;
        END
    END d
END NOR4_Y80

MACRO NOR4_Z1
    CLASS CORE ;
    FOREIGN NOR4_Z1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.090 0.53 1.455 ;
        RECT 0.465 0.090 0.79 0.155 ;
        RECT 0.715 0.090 0.78 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.145 0.530 1.34 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.890 0.530 1.085 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.045 0.530 0.305 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.635 0.530 0.83 0.66 ;
        END
    END d
END NOR4_Z1

MACRO NOR4_Z2
    CLASS CORE ;
    FOREIGN NOR4_Z2 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.040 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.090 1.12 1.455 ;
        RECT 0.925 0.090 1.575 0.155 ;
        RECT 1.425 0.090 1.62 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.285 0.530 2.61 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.780 0.530 2.105 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.085 0.530 0.605 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.275 0.530 1.6 0.66 ;
        END
    END d
END NOR4_Z2

MACRO NOR4_Z3
    CLASS CORE ;
    FOREIGN NOR4_Z3 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 3.800 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.160 0.090 1.355 1.455 ;
        RECT 1.160 0.090 2.005 0.155 ;
        RECT 1.785 0.090 1.98 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.860 0.530 3.25 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.225 0.530 2.615 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.110 0.530 0.76 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.590 0.530 1.98 0.66 ;
        END
    END d
END NOR4_Z3

MACRO NOR4_Z4
    CLASS CORE ;
    FOREIGN NOR4_Z4 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 4.560 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.390 0.090 1.65 1.455 ;
        RECT 1.390 0.090 2.43 0.155 ;
        RECT 2.140 0.090 2.4 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.430 0.530 3.95 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.670 0.530 3.19 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.130 0.530 0.91 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.910 0.530 2.43 0.66 ;
        END
    END d
END NOR4_Z4

MACRO NOR4_Z6
    CLASS CORE ;
    FOREIGN NOR4_Z6 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 5.320 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.620 0.090 1.945 1.455 ;
        RECT 1.620 0.090 2.79 0.155 ;
        RECT 2.495 0.090 2.82 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.000 0.530 4.585 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.115 0.530 3.7 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.150 0.530 1.06 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.230 0.530 2.815 0.66 ;
        END
    END d
END NOR4_Z6

MACRO NOR4_Z8
    CLASS CORE ;
    FOREIGN NOR4_Z8 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.080 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.855 0.090 2.18 1.455 ;
        RECT 1.855 0.090 3.22 0.155 ;
        RECT 2.855 0.090 3.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.575 0.530 5.225 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.560 0.530 4.21 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.175 0.530 1.215 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.545 0.530 3.195 0.66 ;
        END
    END d
END NOR4_Z8

MACRO NOR4_Z10
    CLASS CORE ;
    FOREIGN NOR4_Z10 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 6.460 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 1.970 0.090 2.36 1.455 ;
        RECT 1.970 0.090 3.4 0.155 ;
        RECT 3.030 0.090 3.42 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.860 0.530 5.575 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.785 0.530 4.5 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.185 0.530 1.29 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.705 0.530 3.42 0.66 ;
        END
    END d
END NOR4_Z10

MACRO NOR4_Z20
    CLASS CORE ;
    FOREIGN NOR4_Z20 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 8.740 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 2.665 0.090 3.185 1.455 ;
        RECT 2.665 0.090 4.615 0.155 ;
        RECT 4.100 0.090 4.62 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.575 0.530 7.55 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.115 0.530 6.09 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.250 0.530 1.68 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.660 0.530 4.635 0.66 ;
        END
    END d
END NOR4_Z20

MACRO NOR4_Z40
    CLASS CORE ;
    FOREIGN NOR4_Z40 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 11.780 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 3.590 0.090 4.24 1.455 ;
        RECT 3.590 0.090 6.19 0.155 ;
        RECT 5.530 0.090 6.18 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.860 0.530 10.16 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.895 0.530 8.195 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.335 0.530 2.285 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.935 0.530 6.235 0.66 ;
        END
    END d
END NOR4_Z40

MACRO NOR4_Z80
    CLASS CORE ;
    FOREIGN NOR4_Z80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 16.340 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 4.980 0.090 5.89 1.455 ;
        RECT 4.980 0.090 8.62 0.155 ;
        RECT 7.670 0.090 8.58 0.48 ;
        END
    END o
    PIN a
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 12.290 0.530 14.11 0.66 ;
        END
    END a
    PIN b
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 9.565 0.530 11.385 0.66 ;
        END
    END b
    PIN c
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.465 0.530 3.195 0.66 ;
        END
    END c
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 6.845 0.530 8.665 0.66 ;
        END
    END d
END NOR4_Z80

MACRO DFF_X80
    CLASS CORE ;
    FOREIGN DFF_X80 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 9.500 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN q
        DIRECTION OUTPUT ;
        PORT
        LAYER metal1 ;
        RECT 0.190 0.150 0.45 1.58 ;
        RECT 0.190 0.635 0.775 0.7 ;
        RECT 0.190 1.140 1.62 1.205 ;
        END
    END q
    PIN ck
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 5.240 0.990 5.5 1.38 ;
        RECT 5.240 0.990 5.565 1.185 ;
        RECT 1.815 0.640 2.075 0.835 ;
        RECT 1.565 0.780 2.02 0.845 ;
        RECT 1.815 0.640 3.505 0.705 ;
        RECT 2.815 0.640 3.53 0.835 ;
        RECT 4.330 0.705 4.785 0.835 ;
        RECT 2.815 0.790 4.83 0.855 ;
        RECT 4.580 0.705 4.84 1.03 ;
        RECT 4.580 1.015 5.685 1.08 ;
        RECT 5.190 1.015 5.645 1.145 ;
        RECT 5.240 1.290 5.5 1.485 ;
        RECT 7.940 0.775 8.46 0.84 ;
        RECT 8.240 0.775 8.5 1.49 ;
        RECT 5.240 1.470 8.49 1.535 ;
        RECT 5.240 1.315 5.5 1.38 ;
        RECT 5.315 1.110 5.575 1.175 ;
        RECT 5.315 1.015 5.575 1.08 ;
        END
    END ck
    PIN d
        DIRECTION INPUT ;
        PORT
        LAYER metal1 ;
        RECT 8.705 0.720 8.965 0.785 ;
        END
    END d
END DFF_X80

MACRO TIEH_X1
    CLASS CORE ;
    FOREIGN TIEH_X1 0.000 0.000 ;
    ORIGIN 0.000 0.000 ;
    SIZE 1.520 BY 1.71 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN o
        DIRECTION OUTPUT ;
				USE SIGNAL ;
        PORT
        LAYER metal1 ;
        RECT 0.925 0.150 1.12 1.255 ;
        RECT 0.835 0.150 1.225 0.28 ;
        END
    END o
END TIEH_X1

END LIBRARY
